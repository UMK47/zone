//MAIN_TOP

`define	m1_MIPI_RX0_DPHY_RSTN  reg  [ 0:0]	MIPI_RX0_DPHY_RSTN; wire aMIPI_RX0_DPHY_RSTN = MWE&(MAD==15'h0010); wire [ 0:0]	 bMIPI_RX0_DPHY_RSTN = MDI[0:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_RX0_DPHY_RSTN <= 1'h1; 	else if(aMIPI_RX0_DPHY_RSTN) MIPI_RX0_DPHY_RSTN <= (MBE[0:0] & bMIPI_RX0_DPHY_RSTN) | (~MBE[0:0] & MIPI_RX0_DPHY_RSTN); end  wire [31:0]	wMIPI_RX0_DPHY_RSTN = {32{MAD==15'h0010}} & {31'd0, MIPI_RX0_DPHY_RSTN};
`define	m1_MIPI_RX0_RSTN      reg  [ 0:0]	MIPI_RX0_RSTN; wire aMIPI_RX0_RSTN = MWE&(MAD==15'h0010); wire [ 0:0]	 bMIPI_RX0_RSTN = MDI[1:1]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_RX0_RSTN <= 1'h1; 	else if(aMIPI_RX0_RSTN) MIPI_RX0_RSTN <= (MBE[1:1] & bMIPI_RX0_RSTN) | (~MBE[1:1] & MIPI_RX0_RSTN); end  wire [31:0]	wMIPI_RX0_RSTN = {32{MAD==15'h0010}} & {30'd0, MIPI_RX0_RSTN, 1'd0};
`define	m4_MIPI_RX0_VC_ENA    reg  [ 3:0]	MIPI_RX0_VC_ENA; wire aMIPI_RX0_VC_ENA = MWE&(MAD==15'h0010); wire [ 3:0]	 bMIPI_RX0_VC_ENA = MDI[5:2]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_RX0_VC_ENA <= 4'b0001; 	else if(aMIPI_RX0_VC_ENA) MIPI_RX0_VC_ENA <= (MBE[5:2] & bMIPI_RX0_VC_ENA) | (~MBE[5:2] & MIPI_RX0_VC_ENA); end  wire [31:0]	wMIPI_RX0_VC_ENA = {32{MAD==15'h0010}} & {26'd0, MIPI_RX0_VC_ENA, 2'd0};
`define	m2_MIPI_RX0_LANES     reg  [ 1:0]	MIPI_RX0_LANES; wire aMIPI_RX0_LANES = MWE&(MAD==15'h0010); wire [ 1:0]	 bMIPI_RX0_LANES = MDI[7:6]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_RX0_LANES <= 2'b01; 	else if(aMIPI_RX0_LANES) MIPI_RX0_LANES <= (MBE[7:6] & bMIPI_RX0_LANES) | (~MBE[7:6] & MIPI_RX0_LANES); end  wire [31:0]	wMIPI_RX0_LANES = {32{MAD==15'h0010}} & {24'd0, MIPI_RX0_LANES, 6'd0};
`define	m1_MIPI_RX0_CLEAR     reg  [ 0:0]	MIPI_RX0_CLEAR; wire aMIPI_RX0_CLEAR = MWE&(MAD==15'h0010); wire [ 0:0]	 bMIPI_RX0_CLEAR = MDI[8:8]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_RX0_CLEAR <= 1'h1; 	else if(aMIPI_RX0_CLEAR) MIPI_RX0_CLEAR <= (MBE[8:8] & bMIPI_RX0_CLEAR) | (~MBE[8:8] & MIPI_RX0_CLEAR); end  wire [31:0]	wMIPI_RX0_CLEAR = {32{MAD==15'h0010}} & {23'd0, MIPI_RX0_CLEAR, 8'd0};
`define	m1_MIPI_TX0_DPHY_RSTN  reg  [ 0:0]	MIPI_TX0_DPHY_RSTN; wire aMIPI_TX0_DPHY_RSTN = MWE&(MAD==15'h0011); wire [ 0:0]	 bMIPI_TX0_DPHY_RSTN = MDI[0:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_TX0_DPHY_RSTN <= 1'h1; 	else if(aMIPI_TX0_DPHY_RSTN) MIPI_TX0_DPHY_RSTN <= (MBE[0:0] & bMIPI_TX0_DPHY_RSTN) | (~MBE[0:0] & MIPI_TX0_DPHY_RSTN); end  wire [31:0]	wMIPI_TX0_DPHY_RSTN = {32{MAD==15'h0011}} & {31'd0, MIPI_TX0_DPHY_RSTN};
`define	m1_MIPI_TX0_RSTN      reg  [ 0:0]	MIPI_TX0_RSTN; wire aMIPI_TX0_RSTN = MWE&(MAD==15'h0011); wire [ 0:0]	 bMIPI_TX0_RSTN = MDI[1:1]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_TX0_RSTN <= 1'h1; 	else if(aMIPI_TX0_RSTN) MIPI_TX0_RSTN <= (MBE[1:1] & bMIPI_TX0_RSTN) | (~MBE[1:1] & MIPI_TX0_RSTN); end  wire [31:0]	wMIPI_TX0_RSTN = {32{MAD==15'h0011}} & {30'd0, MIPI_TX0_RSTN, 1'd0};
`define	m2_MIPI_TX0_LANES     reg  [ 1:0]	MIPI_TX0_LANES; wire aMIPI_TX0_LANES = MWE&(MAD==15'h0011); wire [ 1:0]	 bMIPI_TX0_LANES = MDI[3:2]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_TX0_LANES <= 2'b11; 	else if(aMIPI_TX0_LANES) MIPI_TX0_LANES <= (MBE[3:2] & bMIPI_TX0_LANES) | (~MBE[3:2] & MIPI_TX0_LANES); end  wire [31:0]	wMIPI_TX0_LANES = {32{MAD==15'h0011}} & {28'd0, MIPI_TX0_LANES, 2'd0};
`define	m1_MIPI_TX0_FRAME_MODE  reg  [ 0:0]	MIPI_TX0_FRAME_MODE; wire aMIPI_TX0_FRAME_MODE = MWE&(MAD==15'h0011); wire [ 0:0]	 bMIPI_TX0_FRAME_MODE = MDI[7:7]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_TX0_FRAME_MODE <= 1'b0; 	else if(aMIPI_TX0_FRAME_MODE) MIPI_TX0_FRAME_MODE <= (MBE[7:7] & bMIPI_TX0_FRAME_MODE) | (~MBE[7:7] & MIPI_TX0_FRAME_MODE); end  wire [31:0]	wMIPI_TX0_FRAME_MODE = {32{MAD==15'h0011}} & {24'd0, MIPI_TX0_FRAME_MODE, 7'd0};
`define	t16_MIPI_TX0_HRES     reg  [15:0]	_MIPI_TX0_HRES, MIPI_TX0_HRES; wire aMIPI_TX0_HRES = MWE&(MAD==15'h0012); wire [15:0]	 bMIPI_TX0_HRES = MDI[15:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	_MIPI_TX0_HRES <= 16'd1920; 	else if(aMIPI_TX0_HRES) _MIPI_TX0_HRES <= (MBE[15:0] & bMIPI_TX0_HRES) | (~MBE[15:0] & _MIPI_TX0_HRES); end  always @(posedge MTCK or negedge RSTN) begin 	if(!RSTN)	MIPI_TX0_HRES <= 16'd1920; 	else if(VLOCK) MIPI_TX0_HRES <= _MIPI_TX0_HRES; end  wire [31:0]	wMIPI_TX0_HRES = {32{MAD==15'h0012}} & {16'd0, _MIPI_TX0_HRES};
`define	m6_MIPI_TX0_TYPE      reg  [ 5:0]	MIPI_TX0_TYPE; wire aMIPI_TX0_TYPE = MWE&(MAD==15'h0012); wire [ 5:0]	 bMIPI_TX0_TYPE = MDI[21:16]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_TX0_TYPE <= 6'h1e; 	else if(aMIPI_TX0_TYPE) MIPI_TX0_TYPE <= (MBE[21:16] & bMIPI_TX0_TYPE) | (~MBE[21:16] & MIPI_TX0_TYPE); end  wire [31:0]	wMIPI_TX0_TYPE = {32{MAD==15'h0012}} & {10'd0, MIPI_TX0_TYPE, 16'd0};
`define	m2_MIPI_TX0_VC        reg  [ 1:0]	MIPI_TX0_VC; wire aMIPI_TX0_VC = MWE&(MAD==15'h0011); wire [ 1:0]	 bMIPI_TX0_VC = MDI[5:4]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_TX0_VC <= 2'b00; 	else if(aMIPI_TX0_VC) MIPI_TX0_VC <= (MBE[5:4] & bMIPI_TX0_VC) | (~MBE[5:4] & MIPI_TX0_VC); end  wire [31:0]	wMIPI_TX0_VC = {32{MAD==15'h0011}} & {26'd0, MIPI_TX0_VC, 4'd0};
`define	m1_MIPI_TX0_ULPS_CLK_ENTER  reg  [ 0:0]	MIPI_TX0_ULPS_CLK_ENTER; wire aMIPI_TX0_ULPS_CLK_ENTER = MWE&(MAD==15'h0013); wire [ 0:0]	 bMIPI_TX0_ULPS_CLK_ENTER = MDI[0:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_TX0_ULPS_CLK_ENTER <= 1'h0; 	else if(aMIPI_TX0_ULPS_CLK_ENTER) MIPI_TX0_ULPS_CLK_ENTER <= (MBE[0:0] & bMIPI_TX0_ULPS_CLK_ENTER) | (~MBE[0:0] & MIPI_TX0_ULPS_CLK_ENTER); end  wire [31:0]	wMIPI_TX0_ULPS_CLK_ENTER = {32{MAD==15'h0013}} & {31'd0, MIPI_TX0_ULPS_CLK_ENTER};
`define	m1_MIPI_TX0_ULPS_CLK_EXIT  reg  [ 0:0]	MIPI_TX0_ULPS_CLK_EXIT; wire aMIPI_TX0_ULPS_CLK_EXIT = MWE&(MAD==15'h0013); wire [ 0:0]	 bMIPI_TX0_ULPS_CLK_EXIT = MDI[1:1]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_TX0_ULPS_CLK_EXIT <= 1'h0; 	else if(aMIPI_TX0_ULPS_CLK_EXIT) MIPI_TX0_ULPS_CLK_EXIT <= (MBE[1:1] & bMIPI_TX0_ULPS_CLK_EXIT) | (~MBE[1:1] & MIPI_TX0_ULPS_CLK_EXIT); end  wire [31:0]	wMIPI_TX0_ULPS_CLK_EXIT = {32{MAD==15'h0013}} & {30'd0, MIPI_TX0_ULPS_CLK_EXIT, 1'd0};
`define	m4_MIPI_TX0_ULPS_ENTER  reg  [ 3:0]	MIPI_TX0_ULPS_ENTER; wire aMIPI_TX0_ULPS_ENTER = MWE&(MAD==15'h0013); wire [ 3:0]	 bMIPI_TX0_ULPS_ENTER = MDI[7:4]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_TX0_ULPS_ENTER <= 4'h0; 	else if(aMIPI_TX0_ULPS_ENTER) MIPI_TX0_ULPS_ENTER <= (MBE[7:4] & bMIPI_TX0_ULPS_ENTER) | (~MBE[7:4] & MIPI_TX0_ULPS_ENTER); end  wire [31:0]	wMIPI_TX0_ULPS_ENTER = {32{MAD==15'h0013}} & {24'd0, MIPI_TX0_ULPS_ENTER, 4'd0};
`define	m4_MIPI_TX0_ULPS_EXIT  reg  [ 3:0]	MIPI_TX0_ULPS_EXIT; wire aMIPI_TX0_ULPS_EXIT = MWE&(MAD==15'h0013); wire [ 3:0]	 bMIPI_TX0_ULPS_EXIT = MDI[11:8]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MIPI_TX0_ULPS_EXIT <= 4'h0; 	else if(aMIPI_TX0_ULPS_EXIT) MIPI_TX0_ULPS_EXIT <= (MBE[11:8] & bMIPI_TX0_ULPS_EXIT) | (~MBE[11:8] & MIPI_TX0_ULPS_EXIT); end  wire [31:0]	wMIPI_TX0_ULPS_EXIT = {32{MAD==15'h0013}} & {20'd0, MIPI_TX0_ULPS_EXIT, 8'd0};
`define	m1_SS_RSTN            reg  [ 0:0]	SS_RSTN; wire aSS_RSTN = MWE&(MAD==15'h001f); wire [ 0:0]	 bSS_RSTN = MDI[0:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	SS_RSTN <= 1'd1; 	else if(aSS_RSTN) SS_RSTN <= (MBE[0:0] & bSS_RSTN) | (~MBE[0:0] & SS_RSTN); end  wire [31:0]	wSS_RSTN = {32{MAD==15'h001f}} & {31'd0, SS_RSTN};

`define wMAIN_TOP	wire [31:0]	W_MAIN_TOP=wMIPI_RX0_DPHY_RSTN|wMIPI_RX0_RSTN|wMIPI_RX0_VC_ENA|wMIPI_RX0_LANES|wMIPI_RX0_CLEAR|wMIPI_TX0_DPHY_RSTN|wMIPI_TX0_RSTN|wMIPI_TX0_LANES|wMIPI_TX0_FRAME_MODE|wMIPI_TX0_HRES|wMIPI_TX0_TYPE|wMIPI_TX0_VC|wMIPI_TX0_ULPS_CLK_ENTER|wMIPI_TX0_ULPS_CLK_EXIT|wMIPI_TX0_ULPS_ENTER|wMIPI_TX0_ULPS_EXIT|wSS_RSTN;


`define	m6_MIPI_RX0_TYPE       wire [31:0]	rMIPI_RX0_TYPE = {32{MAD==15'h000b}} & {26'd0, MIPI_RX0_TYPE};
`define	m18_MIPI_RX0_ERROR     wire [31:0]	rMIPI_RX0_ERROR = {32{MAD==15'h000c}} & {14'd0, MIPI_RX0_ERROR};
`define	m2_MIPI_RX0_VC         wire [31:0]	rMIPI_RX0_VC = {32{MAD==15'h000b}} & {22'd0, MIPI_RX0_VC, 8'd0};

`define rMAIN_TOP	wire [31:0]	R_MAIN_TOP=rMIPI_RX0_TYPE|rMIPI_RX0_ERROR|rMIPI_RX0_VC;

//SYNC_TOP

`define	m11_SYNC_HSP          reg  [10:0]	SYNC_HSP; wire aSYNC_HSP = MWE&(MAD==15'h0020); wire [10:0]	 bSYNC_HSP = MDI[10:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	SYNC_HSP <= 11'd1; 	else if(aSYNC_HSP) SYNC_HSP <= (MBE[10:0] & bSYNC_HSP) | (~MBE[10:0] & SYNC_HSP); end  wire [31:0]	wSYNC_HSP = {32{MAD==15'h0020}} & {21'd0, SYNC_HSP};
`define	m11_SYNC_VSP          reg  [10:0]	SYNC_VSP; wire aSYNC_VSP = MWE&(MAD==15'h0021); wire [10:0]	 bSYNC_VSP = MDI[10:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	SYNC_VSP <= 11'd28; 	else if(aSYNC_VSP) SYNC_VSP <= (MBE[10:0] & bSYNC_VSP) | (~MBE[10:0] & SYNC_VSP); end  wire [31:0]	wSYNC_VSP = {32{MAD==15'h0021}} & {21'd0, SYNC_VSP};
`define	m12_SYNC_HTW          reg  [11:0]	SYNC_HTW; wire aSYNC_HTW = MWE&(MAD==15'h0016); wire [11:0]	 bSYNC_HTW = MDI[11:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	SYNC_HTW <= 12'd2200; 	else if(aSYNC_HTW) SYNC_HTW <= (MBE[11:0] & bSYNC_HTW) | (~MBE[11:0] & SYNC_HTW); end  wire [31:0]	wSYNC_HTW = {32{MAD==15'h0016}} & {20'd0, SYNC_HTW};
`define	m11_SYNC_VTW          reg  [10:0]	SYNC_VTW; wire aSYNC_VTW = MWE&(MAD==15'h0017); wire [10:0]	 bSYNC_VTW = MDI[10:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	SYNC_VTW <= 11'd1125; 	else if(aSYNC_VTW) SYNC_VTW <= (MBE[10:0] & bSYNC_VTW) | (~MBE[10:0] & SYNC_VTW); end  wire [31:0]	wSYNC_VTW = {32{MAD==15'h0017}} & {21'd0, SYNC_VTW};
`define	m11_SYNC_HW           reg  [10:0]	SYNC_HW; wire aSYNC_HW = MWE&(MAD==15'h0018); wire [10:0]	 bSYNC_HW = MDI[10:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	SYNC_HW <= 11'd1920; 	else if(aSYNC_HW) SYNC_HW <= (MBE[10:0] & bSYNC_HW) | (~MBE[10:0] & SYNC_HW); end  wire [31:0]	wSYNC_HW = {32{MAD==15'h0018}} & {21'd0, SYNC_HW};
`define	m11_SYNC_VW           reg  [10:0]	SYNC_VW; wire aSYNC_VW = MWE&(MAD==15'h0019); wire [10:0]	 bSYNC_VW = MDI[10:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	SYNC_VW <= 11'd1080; 	else if(aSYNC_VW) SYNC_VW <= (MBE[10:0] & bSYNC_VW) | (~MBE[10:0] & SYNC_VW); end  wire [31:0]	wSYNC_VW = {32{MAD==15'h0019}} & {21'd0, SYNC_VW};
`define	m3_CH                 reg  [ 2:0]	CH; wire aCH = MWE&(MAD==15'h002a); wire [ 2:0]	 bCH = MDI[2:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	CH <= 3'd0; 	else if(aCH) CH <= (MBE[2:0] & bCH) | (~MBE[2:0] & CH); end  wire [31:0]	wCH = {32{MAD==15'h002a}} & {29'd0, CH};
`define	m1_SYNC_UP            reg  [ 0:0]	SYNC_UP; wire aSYNC_UP = MWE&(MAD==15'h002b); wire [ 0:0]	 bSYNC_UP = MDI[0:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	SYNC_UP <= 1'd0; 	else if(aSYNC_UP) SYNC_UP <= (MBE[0:0] & bSYNC_UP) | (~MBE[0:0] & SYNC_UP); end  wire [31:0]	wSYNC_UP = {32{MAD==15'h002b}} & {31'd0, SYNC_UP};
`define	m12_DOT_H             reg  [11:0]	DOT_H; wire aDOT_H = MWE&(MAD==15'h0030); wire [11:0]	 bDOT_H = MDI[11:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	DOT_H <= 12'd960; 	else if(aDOT_H) DOT_H <= (MBE[11:0] & bDOT_H) | (~MBE[11:0] & DOT_H); end  wire [31:0]	wDOT_H = {32{MAD==15'h0030}} & {20'd0, DOT_H};
`define	m12_DOT_V             reg  [11:0]	DOT_V; wire aDOT_V = MWE&(MAD==15'h0031); wire [11:0]	 bDOT_V = MDI[11:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	DOT_V <= 12'd540; 	else if(aDOT_V) DOT_V <= (MBE[11:0] & bDOT_V) | (~MBE[11:0] & DOT_V); end  wire [31:0]	wDOT_V = {32{MAD==15'h0031}} & {20'd0, DOT_V};
`define	m12_DOT_W             reg  [11:0]	DOT_W; wire aDOT_W = MWE&(MAD==15'h0032); wire [11:0]	 bDOT_W = MDI[11:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	DOT_W <= 12'd10; 	else if(aDOT_W) DOT_W <= (MBE[11:0] & bDOT_W) | (~MBE[11:0] & DOT_W); end  wire [31:0]	wDOT_W = {32{MAD==15'h0032}} & {20'd0, DOT_W};

`define wSYNC_TOP	wire [31:0]	W_SYNC_TOP=wSYNC_HSP|wSYNC_VSP|wSYNC_HTW|wSYNC_VTW|wSYNC_HW|wSYNC_VW|wCH|wSYNC_UP|wDOT_H|wDOT_V|wDOT_W;

//MTX_TOP

`define	m11_MTX_HTW           reg  [10:0]	MTX_HTW; wire aMTX_HTW = MWE&(MAD==15'h0022); wire [10:0]	 bMTX_HTW = MDI[10:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MTX_HTW <= 11'd1100; 	else if(aMTX_HTW) MTX_HTW <= (MBE[10:0] & bMTX_HTW) | (~MBE[10:0] & MTX_HTW); end  wire [31:0]	wMTX_HTW = {32{MAD==15'h0022}} & {21'd0, MTX_HTW};
`define	m11_MTX_VTW           reg  [10:0]	MTX_VTW; wire aMTX_VTW = MWE&(MAD==15'h0023); wire [10:0]	 bMTX_VTW = MDI[10:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MTX_VTW <= 11'd1125; 	else if(aMTX_VTW) MTX_VTW <= (MBE[10:0] & bMTX_VTW) | (~MBE[10:0] & MTX_VTW); end  wire [31:0]	wMTX_VTW = {32{MAD==15'h0023}} & {21'd0, MTX_VTW};
`define	m11_MTX_HW            reg  [10:0]	MTX_HW; wire aMTX_HW = MWE&(MAD==15'h0024); wire [10:0]	 bMTX_HW = MDI[10:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MTX_HW <= 11'd480; 	else if(aMTX_HW) MTX_HW <= (MBE[10:0] & bMTX_HW) | (~MBE[10:0] & MTX_HW); end  wire [31:0]	wMTX_HW = {32{MAD==15'h0024}} & {21'd0, MTX_HW};
`define	m11_MTX_VW            reg  [10:0]	MTX_VW; wire aMTX_VW = MWE&(MAD==15'h0025); wire [10:0]	 bMTX_VW = MDI[10:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MTX_VW <= 11'd1080; 	else if(aMTX_VW) MTX_VW <= (MBE[10:0] & bMTX_VW) | (~MBE[10:0] & MTX_VW); end  wire [31:0]	wMTX_VW = {32{MAD==15'h0025}} & {21'd0, MTX_VW};
`define	m11_MTX_HSP           reg  [10:0]	MTX_HSP; wire aMTX_HSP = MWE&(MAD==15'h0026); wire [10:0]	 bMTX_HSP = MDI[10:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MTX_HSP <= 11'd481; 	else if(aMTX_HSP) MTX_HSP <= (MBE[10:0] & bMTX_HSP) | (~MBE[10:0] & MTX_HSP); end  wire [31:0]	wMTX_HSP = {32{MAD==15'h0026}} & {21'd0, MTX_HSP};
`define	m11_MTX_VSP           reg  [10:0]	MTX_VSP; wire aMTX_VSP = MWE&(MAD==15'h0027); wire [10:0]	 bMTX_VSP = MDI[10:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MTX_VSP <= 11'd28; 	else if(aMTX_VSP) MTX_VSP <= (MBE[10:0] & bMTX_VSP) | (~MBE[10:0] & MTX_VSP); end  wire [31:0]	wMTX_VSP = {32{MAD==15'h0027}} & {21'd0, MTX_VSP};
`define	m5_HSYNC_WING         reg  [ 4:0]	HSYNC_WING; wire aHSYNC_WING = MWE&(MAD==15'h0028); wire [ 4:0]	 bHSYNC_WING = MDI[9:5]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	HSYNC_WING <= 5'd30; 	else if(aHSYNC_WING) HSYNC_WING <= (MBE[9:5] & bHSYNC_WING) | (~MBE[9:5] & HSYNC_WING); end  wire [31:0]	wHSYNC_WING = {32{MAD==15'h0028}} & {22'd0, HSYNC_WING, 5'd0};
`define	m5_VSYNC_WING         reg  [ 4:0]	VSYNC_WING; wire aVSYNC_WING = MWE&(MAD==15'h0029); wire [ 4:0]	 bVSYNC_WING = MDI[4:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	VSYNC_WING <= 5'd5; 	else if(aVSYNC_WING) VSYNC_WING <= (MBE[4:0] & bVSYNC_WING) | (~MBE[4:0] & VSYNC_WING); end  wire [31:0]	wVSYNC_WING = {32{MAD==15'h0029}} & {27'd0, VSYNC_WING};
`define	t1_MTX_ON             reg  [ 0:0]	_MTX_ON, MTX_ON; wire aMTX_ON = MWE&(MAD==15'h0022); wire [ 0:0]	 bMTX_ON = MDI[31:31]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	_MTX_ON <= 1'd1; 	else if(aMTX_ON) _MTX_ON <= (MBE[31:31] & bMTX_ON) | (~MBE[31:31] & _MTX_ON); end  always @(posedge MTCK or negedge RSTN) begin 	if(!RSTN)	MTX_ON <= 1'd1; 	else if(FLAG_MTCK_RE) MTX_ON <= _MTX_ON; end  wire [31:0]	wMTX_ON = {32{MAD==15'h0022}} & {_MTX_ON, 31'd0};

`define wMTX_TOP	wire [31:0]	W_MTX_TOP=wMTX_HTW|wMTX_VTW|wMTX_HW|wMTX_VW|wMTX_HSP|wMTX_VSP|wHSYNC_WING|wVSYNC_WING|wMTX_ON;

//MRX_TOP

`define	m12_MRX_WR_HW         reg  [11:0]	MRX_WR_HW; wire aMRX_WR_HW = MWE&(MAD==15'h002e); wire [11:0]	 bMRX_WR_HW = MDI[11:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MRX_WR_HW <= 12'd480; 	else if(aMRX_WR_HW) MRX_WR_HW <= (MBE[11:0] & bMRX_WR_HW) | (~MBE[11:0] & MRX_WR_HW); end  wire [31:0]	wMRX_WR_HW = {32{MAD==15'h002e}} & {20'd0, MRX_WR_HW};
`define	m12_MRX_R_HTW         reg  [11:0]	MRX_R_HTW; wire aMRX_R_HTW = MWE&(MAD==15'h002f); wire [11:0]	 bMRX_R_HTW = MDI[11:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MRX_R_HTW <= 12'd2200; 	else if(aMRX_R_HTW) MRX_R_HTW <= (MBE[11:0] & bMRX_R_HTW) | (~MBE[11:0] & MRX_R_HTW); end  wire [31:0]	wMRX_R_HTW = {32{MAD==15'h002f}} & {20'd0, MRX_R_HTW};
`define	m12_MRX_R_VTW         reg  [11:0]	MRX_R_VTW; wire aMRX_R_VTW = MWE&(MAD==15'h003a); wire [11:0]	 bMRX_R_VTW = MDI[11:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MRX_R_VTW <= 12'd1125; 	else if(aMRX_R_VTW) MRX_R_VTW <= (MBE[11:0] & bMRX_R_VTW) | (~MBE[11:0] & MRX_R_VTW); end  wire [31:0]	wMRX_R_VTW = {32{MAD==15'h003a}} & {20'd0, MRX_R_VTW};
`define	m12_MRX_R_HW          reg  [11:0]	MRX_R_HW; wire aMRX_R_HW = MWE&(MAD==15'h003b); wire [11:0]	 bMRX_R_HW = MDI[11:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MRX_R_HW <= 12'd1920; 	else if(aMRX_R_HW) MRX_R_HW <= (MBE[11:0] & bMRX_R_HW) | (~MBE[11:0] & MRX_R_HW); end  wire [31:0]	wMRX_R_HW = {32{MAD==15'h003b}} & {20'd0, MRX_R_HW};
`define	m12_MRX_R_VW          reg  [11:0]	MRX_R_VW; wire aMRX_R_VW = MWE&(MAD==15'h003c); wire [11:0]	 bMRX_R_VW = MDI[11:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MRX_R_VW <= 12'd1080; 	else if(aMRX_R_VW) MRX_R_VW <= (MBE[11:0] & bMRX_R_VW) | (~MBE[11:0] & MRX_R_VW); end  wire [31:0]	wMRX_R_VW = {32{MAD==15'h003c}} & {20'd0, MRX_R_VW};
`define	m12_MRX_R_HSP         reg  [11:0]	MRX_R_HSP; wire aMRX_R_HSP = MWE&(MAD==15'h002c); wire [11:0]	 bMRX_R_HSP = MDI[11:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MRX_R_HSP <= 12'd0; 	else if(aMRX_R_HSP) MRX_R_HSP <= (MBE[11:0] & bMRX_R_HSP) | (~MBE[11:0] & MRX_R_HSP); end  wire [31:0]	wMRX_R_HSP = {32{MAD==15'h002c}} & {20'd0, MRX_R_HSP};
`define	m12_MRX_R_VSP         reg  [11:0]	MRX_R_VSP; wire aMRX_R_VSP = MWE&(MAD==15'h002d); wire [11:0]	 bMRX_R_VSP = MDI[11:0]; always @(posedge MCK or negedge RSTN) begin 	if(!RSTN)	MRX_R_VSP <= 12'd28; 	else if(aMRX_R_VSP) MRX_R_VSP <= (MBE[11:0] & bMRX_R_VSP) | (~MBE[11:0] & MRX_R_VSP); end  wire [31:0]	wMRX_R_VSP = {32{MAD==15'h002d}} & {20'd0, MRX_R_VSP};

`define wMRX_TOP	wire [31:0]	W_MRX_TOP=wMRX_WR_HW|wMRX_R_HTW|wMRX_R_VTW|wMRX_R_HW|wMRX_R_VW|wMRX_R_HSP|wMRX_R_VSP;

